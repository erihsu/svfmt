class testcase extends base_test; /* base class*/
	int a;
	int b;
	function bit funcname();
		return 1'b1;
	endfunction : funcname
endclass : testcase