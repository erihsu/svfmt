program bac;

endprogram

covergroup cg();
	
endgroup : cg